class diffBankAndRowStimulus;

  rand  logic[11:0] row;
  rand  logic[1:0]  bank;

endclass
