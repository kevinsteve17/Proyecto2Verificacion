class sdrcSB;
    int store[$];
    int dir[$];
    int burstLenght[$];
    int ErrCnt;
endclass
