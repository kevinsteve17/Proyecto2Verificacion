class mem_base_object;
    int addr;
    int bl;
    int data[$];
endclass