class sdrcEnv;
    sdrcSB _sb;
    sdrcMon _mon;
    sdrcDrv _drv;
    

    function new (args);
      $$display("Creating SDRC Environment");
            
    endfunction
endclass