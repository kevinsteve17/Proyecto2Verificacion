class stimulus;
  rand  logic[7:0] value;
  //constraint distribution {value dist { 0  := 1 , 1 := 1 }; } 
endclass
