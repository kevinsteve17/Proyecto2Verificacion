class sdrcSB;
    int store[$];
    int dir[$];
    int burstLenght[$];
endclass