class sdrcSB;
    logic [7:0] store[$];
endclass