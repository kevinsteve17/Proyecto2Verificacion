class sdrcSB;
    int store[$]; // need modification to support R/W out of order
    int dir[$];
    int burstLenght[$];
    int ErrCnt;
endclass